module sync_fifo ( 
  // inputs 
  input clk,
  input resetn,
  input [DIN_WIDTH-1:0] data_in ,
  
  // outputs 
 
  ); 
 
endmodule 
