module hello_world ( 
  // inputs 
 
  // outputs 
 
  ); 
 
endmodule 
