module mult_bin #(parameter WIDTH = 4)
  ( 
  // inputs 
  input [WIDTH-1:0] a,
  input [WIDTH-1:0] b,
  // outputs 
  output [2*WIDTH -1:0] y 
  ); 
wire [WIDTH -1 :0] par [WIDTH-1:0] ;
  assign pa
